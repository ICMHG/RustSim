Simple Voltage Divider Circuit
* Basic voltage divider demonstration
* Input: 5V DC source
* Output: Voltage at node 2 should be 2V (due to 1k and 2k resistor ratio)

V1 1 0 DC 5
R1 1 2 1k
R2 2 0 2k

.op
.end 